LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SUMADOR_RESTADOR IS
	PORT(
	NUM1, NUM2 : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	MODO : IN STD_LOGIC;
	NUMR : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
	COUT : OUT STD_LOGIC
	);
	
END SUMADOR_RESTADOR;

ARCHITECTURE BEHAVIOR OF SUMADOR_RESTADOR IS

COMPONENT FULL_ADDER
	PORT(
	A, B, Ci : IN STD_LOGIC;
	Co, S : OUT STD_LOGIC
	);
	
END COMPONENT;

SIGNAL CarryOUt1, CarryOut2, CarryOut3, Xor_1, Xor_2, Xor_3, Xor_4 : STD_LOGIC;

BEGIN

FULLADDER1 : FULL_ADDER PORT MAP (NUM1(0), Xor_1, MODO, CarryOut1, NUMR(0));
FULLADDER2 : FULL_ADDER PORT MAP (NUM1(1), Xor_2, CarryOut1, CarryOut2, NUMR(1));
FULLADDER3 : FULL_ADDER PORT MAP (NUM1(2), Xor_3, CarryOut2, CarryOut3, NUMR(2));
FULLADDER4 : FULL_ADDER PORT MAP (NUM1(3), Xor_4, CarryOut3, COUT, NUMR(3));

Xor_1 <= NUM2(0) XOR MODO;
Xor_2 <= NUM2(1) XOR MODO;
Xor_3 <= NUM2(2) XOR MODO;
Xor_4 <= NUM2(3) XOR MODO;


END BEHAVIOR;